library ieee;
use ieee.std_logic_1164.all;

entity coder is
	port(
		iX : in std_logic_vector(7 downto 0);
		oY : out std_logic_vector(2 downto 0)
	);
end entity;

architecture Behavioral of coder is
	
begin

	
end architecture;